module microcms

pub fn (c Client) content_meta_list<T>(p ListParams) ?T {}
